library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity FluxoDados is
    generic();
    port();
end entity;

architecture of FluxoDados is
    begin

end architecture;